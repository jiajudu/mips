`timescale 1ns / 1ps
module rom(
    input wire Hclock,
    input wire Hreset,
    input wire Hsize,
    input wire Hwrite,
    input wire[31:0] Hwritedata,
    input wire[8:0] Haddress,
    input wire Hselect,
    input wire ready,
    output reg[31:0] Hreaddata,
    output reg Hready,
    output reg Hresponse
);
    reg[31:0] rom[0:127];
    reg[8:0] address;
    always @ (posedge Hclock) begin
        if(Hreset == 1'b0) begin
        end else if(Hselect==1'b1 && ready==1'b1) begin
            address <= Haddress;		
        end
    end
    always @(*) begin
        Hreaddata <= rom[address[8:2]];
        Hresponse <= 1'b0;
        Hready <= 1'b1;
    end
    always @(*) begin
        rom[0] <= 32'h00000000;
        rom[1] <= 32'h10000001;
        rom[2] <= 32'h00000000;
        rom[3] <= 32'h3c10be00;
        rom[4] <= 32'h3c08464c;
        rom[5] <= 32'h3508457f;
        rom[6] <= 32'h240f0000;
        rom[7] <= 32'h020f7821;
        rom[8] <= 32'h8de90000;
        rom[9] <= 32'h8def0004;
        rom[10] <= 32'h000f7c00;
        rom[11] <= 32'h012f4825;
        rom[12] <= 32'h11090003;
        rom[13] <= 32'h00000000;
        rom[14] <= 32'h10000042;
        rom[15] <= 32'h00000000;
        rom[16] <= 32'h240f0038;
        rom[17] <= 32'h020f7821;
        rom[18] <= 32'h8df10000;
        rom[19] <= 32'h8def0004;
        rom[20] <= 32'h000f7c00;
        rom[21] <= 32'h022f8825;
        rom[22] <= 32'h240f0058;
        rom[23] <= 32'h020f7821;
        rom[24] <= 32'h8df20000;
        rom[25] <= 32'h8def0004;
        rom[26] <= 32'h000f7c00;
        rom[27] <= 32'h024f9025;
        rom[28] <= 32'h3252ffff;
        rom[29] <= 32'h240f0030;
        rom[30] <= 32'h020f7821;
        rom[31] <= 32'h8df30000;
        rom[32] <= 32'h8def0004;
        rom[33] <= 32'h000f7c00;
        rom[34] <= 32'h026f9825;
        rom[35] <= 32'h262f0008;
        rom[36] <= 32'h000f7840;
        rom[37] <= 32'h020f7821;
        rom[38] <= 32'h8df40000;
        rom[39] <= 32'h8def0004;
        rom[40] <= 32'h000f7c00;
        rom[41] <= 32'h028fa025;
        rom[42] <= 32'h262f0010;
        rom[43] <= 32'h000f7840;
        rom[44] <= 32'h020f7821;
        rom[45] <= 32'h8df50000;
        rom[46] <= 32'h8def0004;
        rom[47] <= 32'h000f7c00;
        rom[48] <= 32'h02afa825;
        rom[49] <= 32'h262f0004;
        rom[50] <= 32'h000f7840;
        rom[51] <= 32'h020f7821;
        rom[52] <= 32'h8df60000;
        rom[53] <= 32'h8def0004;
        rom[54] <= 32'h000f7c00;
        rom[55] <= 32'h02cfb025;
        rom[56] <= 32'h12800010;
        rom[57] <= 32'h00000000;
        rom[58] <= 32'h12a0000e;
        rom[59] <= 32'h00000000;
        rom[60] <= 32'h26cf0000;
        rom[61] <= 32'h000f7840;
        rom[62] <= 32'h020f7821;
        rom[63] <= 32'h8de80000;
        rom[64] <= 32'h8def0004;
        rom[65] <= 32'h000f7c00;
        rom[66] <= 32'h010f4025;
        rom[67] <= 32'hae880000;
        rom[68] <= 32'h26d60004;
        rom[69] <= 32'h26940004;
        rom[70] <= 32'h26b5fffc;
        rom[71] <= 32'h1ea0fff4;
        rom[72] <= 32'h00000000;
        rom[73] <= 32'h26310020;
        rom[74] <= 32'h2652ffff;
        rom[75] <= 32'h1e40ffd7;
        rom[76] <= 32'h00000000;
        rom[77] <= 32'h02600008;
        rom[78] <= 32'h00000000;
        rom[79] <= 32'h1000ffff;
        rom[80] <= 32'h00000000;
        rom[81] <= 32'h1000ffff;
        rom[82] <= 32'h00000000;
        rom[83] <= 32'h00000000;
        rom[84] <= 32'h00000000;
        rom[85] <= 32'h00000000;
        rom[86] <= 32'h00000000;
        rom[87] <= 32'h00000000;
        rom[88] <= 32'h00000000;
        rom[89] <= 32'h00000000;
        rom[90] <= 32'h00000000;
        rom[91] <= 32'h00000000;
        rom[92] <= 32'h00000000;
        rom[93] <= 32'h00000000;
        rom[94] <= 32'h00000000;
        rom[95] <= 32'h00000000;
        rom[96] <= 32'h00000000;
        rom[97] <= 32'h00000000;
        rom[98] <= 32'h00000000;
        rom[99] <= 32'h00000000;
        rom[100] <= 32'h00000000;
        rom[101] <= 32'h00000000;
        rom[102] <= 32'h00000000;
        rom[103] <= 32'h00000000;
        rom[104] <= 32'h00000000;
        rom[105] <= 32'h00000000;
        rom[106] <= 32'h00000000;
        rom[107] <= 32'h00000000;
        rom[108] <= 32'h00000000;
        rom[109] <= 32'h00000000;
        rom[110] <= 32'h00000000;
        rom[111] <= 32'h00000000;
        rom[112] <= 32'h00000000;
        rom[113] <= 32'h00000000;
        rom[114] <= 32'h00000000;
        rom[115] <= 32'h00000000;
        rom[116] <= 32'h00000000;
        rom[117] <= 32'h00000000;
        rom[118] <= 32'h00000000;
        rom[119] <= 32'h00000000;
        rom[120] <= 32'h00000000;
        rom[121] <= 32'h00000000;
        rom[122] <= 32'h00000000;
        rom[123] <= 32'h00000000;
        rom[124] <= 32'h00000000;
        rom[125] <= 32'h00000000;
        rom[126] <= 32'h00000000;
        rom[127] <= 32'h00000000;
    end
endmodule
