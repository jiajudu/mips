`timescale 1ns / 1ps
module ex_mem(
    input wire clock,
    input wire reset,
    input wire ready,
    input wire flush,
    input wire[31:0] flushTarget,
    input wire[4:0] ExWriteAddress,
    input wire ExWriteRegister,
    input wire[31:0] ExWriteData,
    input wire[31:0] ExWriteHiData,
    input wire[31:0] ExWriteLoData,
    input wire ExWriteHi,
    input wire ExWriteLo,
    input wire ExIsInDelaySlot,
    input wire ExSignExtend,
    input wire ExRAMReadEnable,
    input wire ExWriteCP,
    input wire[4:0] ExWriteCPAddress,
    input wire[31:0] ExWriteCPData,
    input wire Extlbwi,
    input wire Exsyscall,
    input wire Exeret,
    input wire Exprivilege,
    input wire ExValidInstruction,
    input wire PCTLBMiss,
    input wire ExReadTLBMiss,
    input wire ExWriteTLBMiss,
    input wire ExReadError,
    input wire ExWriteError,
    input wire[31:0] ExPC,
    input wire ExAddressReadPrivilege,
    input wire ExAddressWritePrivilege,
    input wire[31:0] ExBadAddress,
    output reg[4:0] MemWriteAddress,
    output reg MemWriteRegister,
    output reg[31:0] MemWriteData,
    output reg[31:0] MemWriteHiData,
    output reg[31:0] MemWriteLoData,
    output reg MemWriteHi,
    output reg MemWriteLo,
    output reg MemIsInDelaySlot,
    output reg MemSignExtend,
    output reg MemRAMReadEnable,
    output reg MemWriteCP,
    output reg[4:0] MemWriteCPAddress,
    output reg[31:0] MemWriteCPData,
    output reg Memtlbwi,
    output reg Memsyscall,
    output reg Memeret,
    output reg Memprivilege,
    output reg TLBMissRead,
    output reg TLBMissWrite,
    output reg ReadError,
    output reg WriteError,
    output reg MemValidInstruction,
    output reg[31:0] MemPC,
    output reg MemAddressReadPrivilege,
    output reg MemAddressWritePrivilege,
    output reg[31:0] MemBadAddress
);
    always @ (posedge clock) begin
        if(reset == 1'b0) begin
            MemWriteAddress <= 5'b00000;
            MemWriteRegister <= 1'b0;
            MemWriteData <= 32'b0;
            MemWriteHiData <= 32'b0;
            MemWriteLoData <= 32'b0;
            MemWriteHi <= 1'b0;
            MemWriteLo <= 1'b0;
            MemRAMReadEnable <= 1'b0;
            MemSignExtend <= 1'b0;
            MemWriteCP <= 1'b0;
            MemWriteCPAddress <= 5'b0;
            MemWriteCPData <= 32'b0;
            Memtlbwi <= 1'b0;
            Memsyscall <= 1'b0;
            Memeret <= 1'b0;
            Memprivilege <= 1'b0;
            MemValidInstruction <= 1'b0;
            TLBMissRead <= 1'b0;
            TLBMissWrite <= 1'b0;
            ReadError <= 1'b0;
            WriteError <= 1'b0;
            MemAddressReadPrivilege <= 1'b0;
            MemAddressWritePrivilege <= 1'b0;
            MemPC <= 32'b0;
            MemBadAddress <= 32'b0;
            MemIsInDelaySlot <= 1'b0;
        end else if(ready == 1'b0) begin
        end else if(flush == 1'b1) begin
            MemWriteAddress <= 5'b00000;
            MemWriteRegister <= 1'b0;
            MemWriteData <= 32'b0;
            MemWriteHiData <= 32'b0;
            MemWriteLoData <= 32'b0;
            MemWriteHi <= 1'b0;
            MemWriteLo <= 1'b0;
            MemRAMReadEnable <= 1'b0;
            MemSignExtend <= 1'b0;
            MemWriteCP <= 1'b0;
            MemWriteCPAddress <= 5'b0;
            MemWriteCPData <= 32'b0;
            Memtlbwi <= 1'b0;
            Memsyscall <= 1'b0;
            Memeret <= 1'b0;
            Memprivilege <= 1'b0;
            MemValidInstruction <= 1'b0;
            TLBMissRead <= 1'b0;
            TLBMissWrite <= 1'b0;
            ReadError <= 1'b0;
            WriteError <= 1'b0;
            MemAddressReadPrivilege <= 1'b0;
            MemAddressWritePrivilege <= 1'b0;
            MemPC <= flushTarget;
            MemBadAddress <= 32'b0;
            MemIsInDelaySlot <= 1'b0;
        end else begin
            MemWriteAddress <= ExWriteAddress;
            MemWriteRegister <= ExWriteRegister;
            MemWriteData <= ExWriteData;
            MemWriteHiData <= ExWriteHiData;
            MemWriteLoData <= ExWriteLoData;
            MemWriteHi <= ExWriteHi;
            MemWriteLo <= ExWriteLo;
            MemRAMReadEnable <= ExRAMReadEnable;
            MemSignExtend <= ExSignExtend;
            MemWriteCP <= ExWriteCP;
            MemWriteCPAddress <= ExWriteCPAddress;
            MemWriteCPData <= ExWriteCPData;
            Memtlbwi <= Extlbwi;
            Memsyscall <= Exsyscall;
            Memeret <= Exeret;
            Memprivilege <= Exprivilege | ExPC[31];
            MemValidInstruction <= ExValidInstruction;
            TLBMissRead <= PCTLBMiss | ExReadTLBMiss;
            TLBMissWrite <= ExWriteTLBMiss;
            ReadError <= ExReadError;
            WriteError <= ExWriteError;
            MemAddressReadPrivilege <= ExAddressReadPrivilege;
            MemAddressWritePrivilege <= ExAddressWritePrivilege;
            MemPC <= ExPC;
            if(PCTLBMiss) begin
                MemBadAddress <= ExPC;
            end else begin
                MemBadAddress <= ExBadAddress;
            end
            MemIsInDelaySlot <= ExIsInDelaySlot;
        end
    end
endmodule