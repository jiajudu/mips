module vga_rom(
    input wire[6:0] ch,
    input wire[6:0] pos,
    output reg mask
);
always @(*) begin
    case(ch[6:0])
        32: begin
            mask = 0;
        end
        33: begin
            case(pos[6:0])
                19, 20, 26, 27, 28, 29, 34, 35, 36, 37, 42, 43, 44, 45, 51, 52, 59, 60, 67, 68, 83, 84, 91, 92:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        34: begin
            case(pos[6:0])
                9, 10, 14, 15, 17, 18, 22, 23, 25, 26, 30, 31, 34, 38:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        35: begin
            case(pos[6:0])
                26, 27, 29, 30, 34, 35, 37, 38, 41, 42, 43, 44, 45, 46, 47, 50, 51, 53, 54, 58, 59, 61, 62, 66, 67, 69, 70, 73, 74, 75, 76, 77, 78, 79, 82, 83, 85, 86, 90, 91, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        36: begin
            case(pos[6:0])
                4, 5, 12, 13, 18, 19, 20, 21, 22, 25, 26, 30, 31, 33, 34, 39, 41, 42, 50, 51, 52, 53, 54, 62, 63, 70, 71, 73, 78, 79, 81, 82, 86, 87, 90, 91, 92, 93, 94, 100, 101, 108, 109:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        37: begin
            case(pos[6:0])
                41, 42, 47, 49, 50, 54, 55, 61, 62, 68, 69, 75, 76, 82, 83, 86, 87, 89, 90, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        38: begin
            case(pos[6:0])
                27, 28, 29, 34, 35, 37, 38, 42, 43, 45, 46, 51, 52, 53, 58, 59, 60, 62, 63, 65, 66, 68, 69, 70, 73, 74, 77, 78, 81, 82, 85, 86, 90, 91, 92, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        39: begin
            case(pos[6:0])
                10, 11, 18, 19, 26, 27, 33, 34:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        40: begin
            case(pos[6:0])
                20, 21, 27, 28, 35, 36, 42, 43, 50, 51, 58, 59, 66, 67, 75, 76, 83, 84, 92, 93:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        41: begin
            case(pos[6:0])
                19, 20, 28, 29, 36, 37, 45, 46, 53, 54, 61, 62, 69, 70, 76, 77, 84, 85, 91, 92:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        42: begin
            case(pos[6:0])
                33, 38, 41, 42, 45, 46, 50, 51, 52, 53, 56, 57, 58, 59, 60, 61, 62, 63, 66, 67, 68, 69, 73, 74, 77, 78, 81, 86:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        43: begin
            case(pos[6:0])
                35, 36, 43, 44, 51, 52, 56, 57, 58, 59, 60, 61, 62, 63, 67, 68, 75, 76, 83, 84:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        44: begin
            case(pos[6:0])
                83, 84, 91, 92, 99, 100, 106, 107:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        45: begin
            case(pos[6:0])
                56, 57, 58, 59, 60, 61, 62, 63:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        46: begin
            case(pos[6:0])
                83, 84, 91, 92:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        47: begin
            case(pos[6:0])
                23, 30, 31, 37, 38, 39, 44, 45, 46, 51, 52, 53, 58, 59, 60, 65, 66, 67, 72, 73, 74, 80, 81, 88:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        48: begin
            case(pos[6:0])
                18, 19, 20, 21, 22, 25, 26, 30, 31, 33, 34, 38, 39, 41, 42, 46, 47, 49, 50, 52, 54, 55, 57, 58, 60, 62, 63, 65, 66, 70, 71, 73, 74, 78, 79, 81, 82, 86, 87, 90, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        49: begin
            case(pos[6:0])
                20, 21, 27, 28, 29, 34, 35, 36, 37, 44, 45, 52, 53, 60, 61, 68, 69, 76, 77, 84, 85, 90, 91, 92, 93, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        50: begin
            case(pos[6:0])
                18, 19, 20, 21, 22, 25, 26, 30, 31, 38, 39, 45, 46, 52, 53, 59, 60, 66, 67, 73, 74, 79, 81, 82, 86, 87, 89, 90, 91, 92, 93, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        51: begin
            case(pos[6:0])
                18, 19, 20, 21, 22, 25, 26, 30, 31, 38, 39, 46, 47, 51, 52, 53, 54, 62, 63, 70, 71, 78, 79, 81, 82, 86, 87, 90, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        52: begin
            case(pos[6:0])
                21, 22, 28, 29, 30, 35, 36, 37, 38, 42, 43, 45, 46, 49, 50, 53, 54, 57, 58, 61, 62, 65, 66, 67, 68, 69, 70, 71, 77, 78, 85, 86, 92, 93, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        53: begin
            case(pos[6:0])
                17, 18, 19, 20, 21, 22, 23, 25, 26, 33, 34, 41, 42, 49, 50, 51, 52, 53, 54, 62, 63, 70, 71, 73, 74, 78, 79, 81, 82, 83, 86, 87, 90, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        54: begin
            case(pos[6:0])
                19, 20, 21, 26, 27, 33, 34, 41, 42, 49, 50, 51, 52, 53, 54, 57, 58, 62, 63, 65, 66, 70, 71, 73, 74, 78, 79, 81, 82, 86, 87, 90, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        55: begin
            case(pos[6:0])
                17, 18, 19, 20, 21, 22, 23, 25, 26, 30, 31, 38, 39, 45, 46, 53, 54, 60, 61, 68, 69, 75, 76, 83, 84, 91, 92:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        56: begin
            case(pos[6:0])
                18, 19, 20, 21, 22, 25, 26, 30, 31, 33, 34, 38, 39, 41, 42, 46, 47, 50, 51, 52, 53, 54, 57, 58, 62, 63, 65, 66, 70, 71, 73, 74, 78, 79, 81, 82, 86, 87, 90, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        57: begin
            case(pos[6:0])
                18, 19, 20, 21, 22, 25, 26, 30, 31, 33, 34, 38, 39, 41, 42, 46, 47, 49, 50, 54, 55, 58, 59, 60, 61, 62, 63, 70, 71, 78, 79, 85, 86, 90, 91, 92, 93:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        58: begin
            case(pos[6:0])
                43, 44, 51, 52, 83, 84, 91, 92:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        59: begin
            case(pos[6:0])
                43, 44, 51, 52, 83, 84, 91, 92, 99, 100, 106, 107:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        60: begin
            case(pos[6:0])
                29, 30, 36, 37, 43, 44, 50, 51, 57, 58, 66, 67, 75, 76, 84, 85, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        61: begin
            case(pos[6:0])
                49, 50, 51, 52, 53, 54, 73, 74, 75, 76, 77, 78:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        62: begin
            case(pos[6:0])
                25, 26, 34, 35, 43, 44, 52, 53, 61, 62, 68, 69, 75, 76, 82, 83, 89, 90:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        63: begin
            case(pos[6:0])
                18, 19, 20, 21, 22, 25, 26, 30, 31, 33, 34, 38, 39, 45, 46, 52, 53, 60, 61, 68, 69, 84, 85, 92, 93:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        64: begin
            case(pos[6:0])
                18, 19, 20, 21, 22, 25, 26, 30, 31, 33, 34, 38, 39, 41, 42, 44, 45, 46, 47, 49, 50, 52, 54, 55, 57, 58, 60, 62, 63, 65, 66, 68, 69, 70, 73, 74, 81, 82, 90, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        65: begin
            case(pos[6:0])
                20, 27, 28, 29, 34, 35, 37, 38, 41, 42, 46, 47, 49, 50, 54, 55, 57, 58, 62, 63, 65, 66, 67, 68, 69, 70, 71, 73, 74, 78, 79, 81, 82, 86, 87, 89, 90, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        66: begin
            case(pos[6:0])
                17, 18, 19, 20, 21, 22, 26, 27, 30, 31, 34, 35, 38, 39, 42, 43, 46, 47, 50, 51, 52, 53, 54, 58, 59, 62, 63, 66, 67, 70, 71, 74, 75, 78, 79, 82, 83, 86, 87, 89, 90, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        67: begin
            case(pos[6:0])
                19, 20, 21, 22, 26, 27, 30, 31, 33, 34, 39, 41, 42, 49, 50, 57, 58, 65, 66, 73, 74, 79, 82, 83, 86, 87, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        68: begin
            case(pos[6:0])
                17, 18, 19, 20, 21, 26, 27, 29, 30, 34, 35, 38, 39, 42, 43, 46, 47, 50, 51, 54, 55, 58, 59, 62, 63, 66, 67, 70, 71, 74, 75, 78, 79, 82, 83, 85, 86, 89, 90, 91, 92, 93:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        69: begin
            case(pos[6:0])
                17, 18, 19, 20, 21, 22, 23, 26, 27, 30, 31, 34, 35, 39, 42, 43, 45, 50, 51, 52, 53, 58, 59, 61, 66, 67, 74, 75, 79, 82, 83, 86, 87, 89, 90, 91, 92, 93, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        70: begin
            case(pos[6:0])
                17, 18, 19, 20, 21, 22, 23, 26, 27, 30, 31, 34, 35, 39, 42, 43, 45, 50, 51, 52, 53, 58, 59, 61, 66, 67, 74, 75, 82, 83, 89, 90, 91, 92:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        71: begin
            case(pos[6:0])
                19, 20, 21, 22, 26, 27, 30, 31, 33, 34, 39, 41, 42, 49, 50, 57, 58, 60, 61, 62, 63, 65, 66, 70, 71, 73, 74, 78, 79, 82, 83, 85, 86, 87, 91, 92, 93, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        72: begin
            case(pos[6:0])
                17, 18, 22, 23, 25, 26, 30, 31, 33, 34, 38, 39, 41, 42, 46, 47, 49, 50, 51, 52, 53, 54, 55, 57, 58, 62, 63, 65, 66, 70, 71, 73, 74, 78, 79, 81, 82, 86, 87, 89, 90, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        73: begin
            case(pos[6:0])
                18, 19, 20, 21, 27, 28, 35, 36, 43, 44, 51, 52, 59, 60, 67, 68, 75, 76, 83, 84, 90, 91, 92, 93:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        74: begin
            case(pos[6:0])
                20, 21, 22, 23, 29, 30, 37, 38, 45, 46, 53, 54, 61, 62, 69, 70, 73, 74, 77, 78, 81, 82, 85, 86, 90, 91, 92, 93:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        75: begin
            case(pos[6:0])
                17, 18, 19, 22, 23, 26, 27, 30, 31, 34, 35, 37, 38, 42, 43, 45, 46, 50, 51, 52, 53, 58, 59, 61, 62, 66, 67, 69, 70, 74, 75, 78, 79, 82, 83, 86, 87, 89, 90, 91, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        76: begin
            case(pos[6:0])
                17, 18, 19, 20, 26, 27, 34, 35, 42, 43, 50, 51, 58, 59, 66, 67, 74, 75, 79, 82, 83, 86, 87, 89, 90, 91, 92, 93, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        77: begin
            case(pos[6:0])
                17, 18, 22, 23, 25, 26, 27, 29, 30, 31, 33, 34, 35, 36, 37, 38, 39, 41, 42, 44, 46, 47, 49, 50, 54, 55, 57, 58, 62, 63, 65, 66, 70, 71, 73, 74, 78, 79, 81, 82, 86, 87, 89, 90, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        78: begin
            case(pos[6:0])
                17, 18, 22, 23, 25, 26, 30, 31, 33, 34, 35, 38, 39, 41, 42, 43, 44, 46, 47, 49, 50, 51, 52, 53, 54, 55, 57, 58, 60, 61, 62, 63, 65, 66, 69, 70, 71, 73, 74, 78, 79, 81, 82, 86, 87, 89, 90, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        79: begin
            case(pos[6:0])
                19, 20, 21, 26, 27, 29, 30, 33, 34, 38, 39, 41, 42, 46, 47, 49, 50, 54, 55, 57, 58, 62, 63, 65, 66, 70, 71, 73, 74, 78, 79, 82, 83, 85, 86, 91, 92, 93:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        80: begin
            case(pos[6:0])
                17, 18, 19, 20, 21, 22, 26, 27, 30, 31, 34, 35, 38, 39, 42, 43, 46, 47, 50, 51, 52, 53, 54, 58, 59, 66, 67, 74, 75, 82, 83, 89, 90, 91, 92:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        81: begin
            case(pos[6:0])
                18, 19, 20, 21, 22, 25, 26, 30, 31, 33, 34, 38, 39, 41, 42, 46, 47, 49, 50, 54, 55, 57, 58, 62, 63, 65, 66, 70, 71, 73, 74, 76, 78, 79, 81, 82, 84, 85, 86, 87, 90, 91, 92, 93, 94, 101, 102, 109, 110, 111:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        82: begin
            case(pos[6:0])
                17, 18, 19, 20, 21, 22, 26, 27, 30, 31, 34, 35, 38, 39, 42, 43, 46, 47, 50, 51, 52, 53, 54, 58, 59, 61, 62, 66, 67, 69, 70, 74, 75, 78, 79, 82, 83, 86, 87, 89, 90, 91, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        83: begin
            case(pos[6:0])
                18, 19, 20, 21, 22, 25, 26, 30, 31, 33, 34, 38, 39, 42, 43, 51, 52, 53, 61, 62, 70, 71, 73, 74, 78, 79, 81, 82, 86, 87, 90, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        84: begin
            case(pos[6:0])
                16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 27, 28, 30, 31, 32, 35, 36, 39, 43, 44, 51, 52, 59, 60, 67, 68, 75, 76, 83, 84, 90, 91, 92, 93:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        85: begin
            case(pos[6:0])
                17, 18, 22, 23, 25, 26, 30, 31, 33, 34, 38, 39, 41, 42, 46, 47, 49, 50, 54, 55, 57, 58, 62, 63, 65, 66, 70, 71, 73, 74, 78, 79, 81, 82, 86, 87, 90, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        86: begin
            case(pos[6:0])
                17, 18, 22, 23, 25, 26, 30, 31, 33, 34, 38, 39, 41, 42, 46, 47, 49, 50, 54, 55, 57, 58, 62, 63, 65, 66, 70, 71, 74, 75, 77, 78, 83, 84, 85, 92:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        87: begin
            case(pos[6:0])
                17, 18, 22, 23, 25, 26, 30, 31, 33, 34, 38, 39, 41, 42, 46, 47, 49, 50, 54, 55, 57, 58, 60, 62, 63, 65, 66, 68, 70, 71, 73, 74, 75, 76, 77, 78, 79, 82, 83, 85, 86, 90, 91, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        88: begin
            case(pos[6:0])
                16, 17, 22, 23, 24, 25, 30, 31, 33, 34, 37, 38, 42, 43, 44, 45, 51, 52, 59, 60, 66, 67, 68, 69, 73, 74, 77, 78, 80, 81, 86, 87, 88, 89, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        89: begin
            case(pos[6:0])
                16, 17, 22, 23, 24, 25, 30, 31, 32, 33, 38, 39, 41, 42, 45, 46, 50, 51, 52, 53, 59, 60, 67, 68, 75, 76, 83, 84, 90, 91, 92, 93:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        90: begin
            case(pos[6:0])
                17, 18, 19, 20, 21, 22, 23, 25, 26, 30, 31, 33, 38, 39, 45, 46, 52, 53, 59, 60, 66, 67, 73, 74, 79, 81, 82, 86, 87, 89, 90, 91, 92, 93, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        91: begin
            case(pos[6:0])
                18, 19, 20, 21, 26, 27, 34, 35, 42, 43, 50, 51, 58, 59, 66, 67, 74, 75, 82, 83, 90, 91, 92, 93:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        92: begin
            case(pos[6:0])
                16, 24, 25, 32, 33, 34, 41, 42, 43, 50, 51, 52, 59, 60, 61, 68, 69, 70, 77, 78, 79, 86, 87, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        93: begin
            case(pos[6:0])
                18, 19, 20, 21, 28, 29, 36, 37, 44, 45, 52, 53, 60, 61, 68, 69, 76, 77, 84, 85, 90, 91, 92, 93:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        94: begin
            case(pos[6:0])
                4, 11, 12, 13, 18, 19, 21, 22, 25, 26, 30, 31:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        95: begin
            case(pos[6:0])
                96, 97, 98, 99, 100, 101, 102, 103:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        96: begin
            case(pos[6:0])
                3, 4, 11, 12, 20, 21:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        97: begin
            case(pos[6:0])
                42, 43, 44, 45, 49, 53, 54, 61, 62, 66, 67, 68, 69, 70, 73, 74, 77, 78, 81, 82, 85, 86, 90, 91, 92, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        98: begin
            case(pos[6:0])
                17, 18, 19, 26, 27, 34, 35, 42, 43, 44, 45, 50, 51, 53, 54, 58, 59, 62, 63, 66, 67, 70, 71, 74, 75, 78, 79, 82, 83, 86, 87, 89, 90, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        99: begin
            case(pos[6:0])
                42, 43, 44, 45, 46, 49, 50, 54, 55, 57, 58, 65, 66, 73, 74, 81, 82, 86, 87, 90, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        100: begin
            case(pos[6:0])
                20, 21, 22, 29, 30, 37, 38, 43, 44, 45, 46, 50, 51, 53, 54, 57, 58, 61, 62, 65, 66, 69, 70, 73, 74, 77, 78, 81, 82, 85, 86, 90, 91, 92, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        101: begin
            case(pos[6:0])
                42, 43, 44, 45, 46, 49, 50, 54, 55, 57, 58, 62, 63, 65, 66, 67, 68, 69, 70, 73, 74, 81, 82, 86, 87, 90, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        102: begin
            case(pos[6:0])
                19, 20, 21, 26, 27, 29, 30, 34, 35, 38, 42, 43, 49, 50, 51, 52, 53, 58, 59, 66, 67, 74, 75, 82, 83, 89, 90, 91, 92:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        103: begin
            case(pos[6:0])
                42, 43, 44, 46, 47, 49, 50, 53, 54, 57, 58, 61, 62, 65, 66, 69, 70, 73, 74, 77, 78, 82, 83, 84, 85, 86, 93, 94, 97, 98, 101, 102, 106, 107, 108, 109:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        104: begin
            case(pos[6:0])
                17, 18, 19, 26, 27, 34, 35, 42, 43, 45, 46, 50, 51, 52, 54, 55, 58, 59, 62, 63, 66, 67, 70, 71, 74, 75, 78, 79, 82, 83, 86, 87, 89, 90, 91, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        105: begin
            case(pos[6:0])
                20, 21, 28, 29, 43, 44, 45, 52, 53, 60, 61, 68, 69, 76, 77, 84, 85, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        106: begin
            case(pos[6:0])
                21, 22, 29, 30, 44, 45, 46, 53, 54, 61, 62, 69, 70, 77, 78, 85, 86, 89, 90, 93, 94, 97, 98, 101, 102, 106, 107, 108, 109:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        107: begin
            case(pos[6:0])
                17, 18, 19, 26, 27, 34, 35, 42, 43, 46, 47, 50, 51, 54, 55, 58, 59, 61, 62, 66, 67, 68, 69, 74, 75, 77, 78, 82, 83, 86, 87, 89, 90, 91, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        108: begin
            case(pos[6:0])
                19, 20, 21, 28, 29, 36, 37, 44, 45, 52, 53, 60, 61, 68, 69, 76, 77, 84, 85, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        109: begin
            case(pos[6:0])
                41, 42, 44, 45, 46, 49, 50, 51, 52, 53, 54, 55, 57, 58, 60, 62, 63, 65, 66, 68, 70, 71, 73, 74, 76, 78, 79, 81, 82, 84, 86, 87, 89, 90, 92, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        110: begin
            case(pos[6:0])
                41, 42, 44, 45, 46, 50, 51, 54, 55, 58, 59, 62, 63, 66, 67, 70, 71, 74, 75, 78, 79, 82, 83, 86, 87, 90, 91, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        111: begin
            case(pos[6:0])
                42, 43, 44, 45, 46, 49, 50, 54, 55, 57, 58, 62, 63, 65, 66, 70, 71, 73, 74, 78, 79, 81, 82, 86, 87, 90, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        112: begin
            case(pos[6:0])
                41, 42, 44, 45, 46, 50, 51, 54, 55, 58, 59, 62, 63, 66, 67, 70, 71, 74, 75, 78, 79, 82, 83, 84, 85, 86, 90, 91, 98, 99, 105, 106, 107, 108:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        113: begin
            case(pos[6:0])
                42, 43, 44, 46, 47, 49, 50, 53, 54, 57, 58, 61, 62, 65, 66, 69, 70, 73, 74, 77, 78, 82, 83, 84, 85, 86, 93, 94, 101, 102, 108, 109, 110, 111:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        114: begin
            case(pos[6:0])
                41, 42, 44, 45, 46, 50, 51, 52, 54, 55, 58, 59, 62, 63, 66, 67, 74, 75, 82, 83, 89, 90, 91, 92:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        115: begin
            case(pos[6:0])
                42, 43, 44, 45, 46, 49, 50, 54, 55, 58, 59, 60, 68, 69, 70, 78, 79, 81, 82, 86, 87, 90, 91, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        116: begin
            case(pos[6:0])
                20, 27, 28, 35, 36, 41, 42, 43, 44, 45, 46, 51, 52, 59, 60, 67, 68, 75, 76, 83, 84, 86, 87, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        117: begin
            case(pos[6:0])
                41, 42, 45, 46, 49, 50, 53, 54, 57, 58, 61, 62, 65, 66, 69, 70, 73, 74, 77, 78, 81, 82, 85, 86, 90, 91, 92, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        118: begin
            case(pos[6:0])
                41, 42, 46, 47, 49, 50, 54, 55, 58, 59, 61, 62, 66, 67, 69, 70, 75, 76, 77, 83, 84, 85, 92:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        119: begin
            case(pos[6:0])
                41, 42, 46, 47, 49, 50, 54, 55, 57, 58, 62, 63, 65, 66, 68, 70, 71, 73, 74, 76, 78, 79, 81, 82, 83, 84, 85, 86, 87, 90, 91, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        120: begin
            case(pos[6:0])
                41, 42, 46, 47, 50, 51, 53, 54, 59, 60, 61, 67, 68, 69, 75, 76, 77, 82, 83, 85, 86, 89, 90, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        121: begin
            case(pos[6:0])
                41, 42, 46, 47, 49, 50, 54, 55, 57, 58, 62, 63, 65, 66, 70, 71, 73, 74, 78, 79, 82, 83, 84, 85, 86, 87, 94, 95, 101, 102, 106, 107, 108, 109:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        122: begin
            case(pos[6:0])
                41, 42, 43, 44, 45, 46, 47, 49, 50, 53, 54, 60, 61, 67, 68, 74, 75, 81, 82, 86, 87, 89, 90, 91, 92, 93, 94, 95:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        123: begin
            case(pos[6:0])
                20, 21, 22, 27, 28, 35, 36, 43, 44, 49, 50, 51, 59, 60, 67, 68, 75, 76, 83, 84, 92, 93, 94:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        124: begin
            case(pos[6:0])
                19, 20, 27, 28, 35, 36, 43, 44, 51, 52, 67, 68, 75, 76, 83, 84, 91, 92, 99, 100:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        125: begin
            case(pos[6:0])
                17, 18, 19, 27, 28, 35, 36, 43, 44, 52, 53, 54, 59, 60, 67, 68, 75, 76, 83, 84, 89, 90, 91:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        126: begin
            case(pos[6:0])
                18, 19, 20, 22, 23, 25, 26, 28, 29, 30:
                    mask = 1;
                default: mask = 0;
            endcase
        end
        default: begin
            mask = 0;
        end
    endcase
end

endmodule